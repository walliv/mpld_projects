----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
----------------------------------------------------------------------------------
ENTITY FIR_50k_SIM IS
  PORT (
    aclk                                : IN  STD_LOGIC;
    s_axis_data_tvalid                  : IN  STD_LOGIC;
    s_axis_data_tready                  : OUT STD_LOGIC;
    s_axis_data_tdata                   : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
    m_axis_data_tvalid                  : OUT STD_LOGIC := '0';
    m_axis_data_tdata                   : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0')
  );
END FIR_50k_SIM;
----------------------------------------------------------------------------------
ARCHITECTURE structural OF FIR_50k_SIM IS
----------------------------------------------------------------------------------

  SIGNAL cnt_fir_out                    : INTEGER := 0;
  SIGNAL cnt_fir_in                     : INTEGER := 0;
  SIGNAL s_axis_data_tvalid_i           : STD_LOGIC := '0';
  SIGNAL s_axis_data_tvalid_ii          : STD_LOGIC := '0';

  TYPE t_fir_response IS ARRAY (0 TO 999) OF INTEGER;
  CONSTANT C_FIR_RESPONSE               : t_fir_response := (
0,
0,
-1,
-1,
-1,
0,
0,
1,
1,
2,
3,
4,
5,
7,
8,
10,
12,
14,
17,
20,
23,
26,
29,
33,
37,
41,
45,
49,
53,
57,
63,
67,
72,
76,
81,
85,
90,
94,
98,
102,
106,
110,
115,
117,
120,
124,
127,
130,
132,
134,
136,
138,
139,
141,
142,
144,
145,
145,
146,
148,
149,
148,
148,
149,
149,
149,
150,
149,
149,
148,
148,
146,
145,
143,
140,
139,
136,
133,
130,
125,
120,
116,
111,
107,
100,
94,
88,
82,
75,
68,
60,
53,
46,
39,
31,
24,
17,
9,
2,
-5,
-12,
-18,
-24,
-31,
-36,
-42,
-45,
-51,
-55,
-59,
-63,
-67,
-69,
-72,
-73,
-76,
-77,
-80,
-81,
-81,
-83,
-84,
-85,
-84,
-85,
-85,
-85,
-87,
-87,
-87,
-86,
-86,
-84,
-85,
-83,
-82,
-80,
-77,
-76,
-72,
-70,
-66,
-60,
-57,
-52,
-46,
-41,
-33,
-28,
-21,
-13,
-7,
3,
9,
17,
27,
34,
42,
50,
58,
67,
74,
82,
89,
96,
103,
108,
114,
120,
124,
129,
131,
135,
140,
141,
145,
145,
147,
148,
149,
149,
149,
149,
149,
149,
150,
147,
146,
145,
146,
145,
146,
143,
143,
141,
138,
138,
136,
134,
131,
129,
126,
122,
119,
116,
111,
106,
101,
96,
91,
84,
79,
72,
65,
59,
51,
44,
36,
29,
23,
14,
9,
2,
-6,
-12,
-19,
-24,
-29,
-36,
-40,
-46,
-50,
-54,
-59,
-62,
-66,
-69,
-71,
-74,
-75,
-78,
-80,
-81,
-83,
-83,
-85,
-86,
-88,
-88,
-89,
-88,
-89,
-92,
-91,
-91,
-92,
-91,
-91,
-90,
-89,
-87,
-87,
-83,
-80,
-79,
-75,
-71,
-66,
-62,
-57,
-52,
-46,
-38,
-32,
-25,
-18,
-10,
-3,
5,
12,
21,
29,
36,
44,
51,
59,
67,
73,
79,
86,
92,
98,
103,
108,
113,
116,
122,
123,
129,
132,
133,
135,
137,
140,
141,
142,
144,
143,
144,
146,
146,
144,
145,
144,
146,
144,
143,
142,
141,
141,
137,
135,
133,
130,
126,
122,
119,
114,
109,
104,
98,
93,
85,
78,
71,
65,
57,
49,
40,
32,
23,
14,
6,
-3,
-10,
-18,
-27,
-36,
-42,
-50,
-57,
-64,
-70,
-75,
-80,
-85,
-91,
-93,
-96,
-99,
-104,
-107,
-107,
-109,
-111,
-111,
-112,
-114,
-113,
-113,
-113,
-112,
-113,
-110,
-110,
-110,
-109,
-110,
-108,
-107,
-106,
-105,
-103,
-102,
-100,
-98,
-96,
-93,
-90,
-86,
-83,
-79,
-74,
-69,
-63,
-57,
-52,
-46,
-38,
-31,
-23,
-15,
-6,
2,
11,
19,
28,
38,
46,
54,
64,
71,
80,
89,
95,
103,
109,
115,
122,
127,
132,
135,
140,
144,
146,
150,
151,
153,
156,
155,
157,
156,
157,
157,
157,
158,
156,
156,
155,
156,
157,
155,
153,
154,
152,
150,
150,
147,
146,
143,
141,
138,
133,
131,
125,
121,
116,
110,
104,
97,
91,
85,
76,
71,
61,
52,
44,
35,
27,
18,
8,
0,
-8,
-16,
-24,
-33,
-41,
-47,
-53,
-59,
-66,
-70,
-74,
-80,
-83,
-88,
-90,
-91,
-94,
-95,
-97,
-98,
-98,
-99,
-99,
-99,
-98,
-99,
-97,
-95,
-95,
-95,
-95,
-94,
-93,
-92,
-92,
-89,
-89,
-86,
-85,
-83,
-79,
-77,
-73,
-69,
-66,
-61,
-56,
-51,
-46,
-41,
-33,
-25,
-20,
-12,
-5,
3,
10,
18,
27,
34,
43,
50,
57,
64,
72,
79,
86,
90,
96,
102,
107,
112,
114,
118,
122,
123,
126,
127,
129,
131,
130,
132,
131,
132,
131,
131,
131,
131,
131,
128,
127,
127,
128,
127,
127,
125,
125,
123,
122,
121,
119,
118,
117,
112,
110,
107,
103,
99,
94,
89,
85,
79,
74,
67,
61,
54,
47,
40,
32,
25,
17,
8,
0,
-5,
-15,
-20,
-30,
-36,
-44,
-50,
-55,
-63,
-68,
-72,
-78,
-83,
-88,
-92,
-95,
-98,
-101,
-105,
-106,
-110,
-111,
-112,
-113,
-115,
-118,
-119,
-120,
-118,
-118,
-119,
-120,
-121,
-122,
-122,
-120,
-120,
-120,
-119,
-119,
-116,
-115,
-113,
-111,
-108,
-105,
-101,
-97,
-93,
-87,
-82,
-77,
-70,
-66,
-59,
-52,
-44,
-38,
-32,
-23,
-16,
-7,
0,
7,
16,
22,
30,
37,
45,
52,
59,
66,
71,
76,
82,
87,
91,
95,
100,
103,
106,
110,
114,
115,
117,
118,
120,
124,
124,
125,
126,
126,
126,
125,
129,
129,
129,
127,
127,
128,
126,
124,
123,
120,
119,
116,
114,
111,
107,
105,
98,
95,
90,
84,
77,
73,
66,
59,
51,
45,
37,
29,
22,
15,
5,
-2,
-10,
-18,
-26,
-33,
-40,
-47,
-54,
-60,
-67,
-73,
-77,
-83,
-88,
-93,
-98,
-99,
-103,
-105,
-110,
-111,
-112,
-115,
-116,
-116,
-117,
-118,
-121,
-119,
-119,
-119,
-119,
-121,
-119,
-118,
-118,
-116,
-116,
-115,
-112,
-109,
-106,
-105,
-101,
-98,
-94,
-89,
-83,
-79,
-73,
-68,
-61,
-55,
-46,
-39,
-32,
-24,
-15,
-7,
1,
10,
19,
27,
37,
44,
53,
61,
70,
77,
83,
92,
98,
104,
109,
114,
120,
125,
129,
132,
135,
138,
140,
142,
144,
144,
146,
147,
146,
147,
146,
147,
144,
144,
143,
144,
143,
141,
139,
138,
137,
135,
132,
129,
126,
124,
120,
116,
112,
107,
104,
98,
92,
88,
80,
75,
67,
61,
55,
47,
40,
30,
23,
16,
9,
-1,
-9,
-16,
-24,
-31,
-38,
-45,
-52,
-59,
-64,
-69,
-74,
-81,
-85,
-90,
-92,
-97,
-100,
-102,
-106,
-108,
-108,
-110,
-111,
-112,
-113,
-114,
-114,
-114,
-113,
-113,
-113,
-112,
-114,
-111,
-111,
-111,
-110,
-109,
-107,
-105,
-103,
-101,
-100,
-96,
-93,
-90,
-85,
-83,
-79,
-74,
-69,
-64,
-59,
-53,
-48,
-43,
-36,
-29,
-24,
-16,
-10,
-5,
2,
8,
15,
22,
27,
34,
40,
46,
52,
57,
60,
66,
70,
75,
80,
83,
86,
91,
94,
96,
100,
101,
104,
107,
109,
110,
113,
114,
117,
115,
118,
119,
122,
122,
123,
123,
123,
124,
124,
122,
122,
120,
119,
118,
115,
112,
109,
105,
101,
96,
92,
87,
80,
75,
67,
61,
55,
47,
39,
31,
24,
16,
8,
0,
-6,
-14,
-21,
-28,
-34,
-40,
-48,
-53,
-58,
-64,
-69,
-74,
-76,
-80,
-84,
-85,
-89,
-91,
-91,
-92,
-94,
-95,
-94,
-94,
-95,
-95,
-95,
-93,
-93
  );


  CONSTANT C_FIR_IN : t_fir_response := (
127,
128,
127,
127,
193,
127,
143,
131,
131,
160,
136,
127,
127,
209,
127,
147,
163,
132,
160,
200,
193,
143,
65,
127,
144,
131,
131,
226,
136,
143,
131,
213,
160,
156,
163,
132,
242,
200,
213,
179,
70,
160,
215,
197,
147,
32,
136,
128,
127,
209,
193,
147,
179,
128,
164,
231,
202,
143,
65,
209,
144,
143,
-96,
-26,
-88,
-39,
-58,
-58,
-157,
-99,
-75,
-127,
-9,
-86,
-33,
-92,
-189,
-9,
-7,
-37,
-80,
-220,
-6,
-56,
-42,
-26,
-251,
-75,
-20,
-57,
-79,
-183,
-62,
-111,
-190,
-128,
-45,
-124,
-108,
-25,
-115,
-79,
-115,
-42,
-95,
-49,
-92,
-111,
-41,
-52,
-9,
-3,
-251,
-79,
-230,
-58,
-123,
-219,
-115,
-30,
-119,
-62,
-58,
-62,
-107,
155,
128,
236,
183,
216,
19,
229,
85,
176,
247,
159,
187,
119,
206,
198,
98,
206,
246,
148,
194,
170,
249,
203,
7,
230,
58,
136,
160,
51,
217,
173,
253,
190,
66,
242,
14,
217,
131,
71,
180,
186,
28,
163,
15,
242,
236,
187,
188,
20,
246,
157,
246,
168,
32,
163,
186,
138,
197,
51,
70,
159,
215,
-58,
-42,
-223,
-103,
-123,
-124,
-13,
-53,
-108,
-76,
-45,
-91,
-4,
-17,
-107,
-157,
-101,
-45,
-128,
-158,
-26,
-71,
-35,
-62,
-91,
-150,
-115,
-79,
-41,
-42,
-73,
-5,
-95,
-208,
-66,
-81,
-17,
-137,
-251,
-94,
-114,
-62,
-185,
-244,
-76,
-20,
-107,
-13,
-163,
-10,
-112,
-153,
-24,
-104,
-108,
-170,
-75,
-100,
-95,
-83,
-80,
-119,
-106,
225,
214,
51,
208,
193,
251,
113,
154,
68,
225,
69,
81,
243,
184,
184,
101,
187,
137,
194,
249,
3,
215,
211,
157,
36,
46,
19,
159,
57,
159,
238,
123,
218,
159,
109,
253,
249,
194,
225,
227,
221,
220,
94,
170,
75,
243,
35,
4,
63,
231,
250,
25,
77,
144,
5,
151,
193,
9,
159,
166,
27,
200,
-216,
-86,
-135,
-38,
-149,
-220,
-113,
-66,
-53,
-175,
-146,
-29,
-168,
-60,
-79,
-223,
-252,
-117,
-94,
-118,
-162,
-186,
-222,
-116,
-91,
-185,
-111,
-70,
-54,
-20,
-154,
-113,
-160,
-49,
-153,
-173,
-26,
-69,
-1,
-62,
-215,
-82,
-81,
-103,
-169,
-232,
-58,
-55,
-95,
-98,
-166,
-123,
-245,
-75,
-23,
-165,
-80,
-219,
-6,
-56,
-108,
-26,
-235,
176,
231,
229,
183,
72,
193,
194,
65,
147,
246,
128,
180,
173,
206,
160,
78,
213,
175,
202,
159,
241,
221,
219,
242,
170,
35,
171,
61,
194,
245,
107,
218,
213,
77,
226,
157,
131,
128,
60,
135,
235,
183,
138,
85,
241,
97,
175,
220,
199,
246,
103,
12,
148,
113,
222,
214,
242,
234,
241,
187,
137,
234,
-6,
-242,
-120,
-42,
-226,
-123,
-118,
-195,
-56,
-198,
-88,
-193,
-130,
-2,
-256,
-29,
-35,
-104,
-111,
-132,
-76,
-36,
-139,
-1,
-252,
-203,
-98,
-92,
-83,
-203,
-61,
-74,
-70,
-53,
-158,
-154,
-17,
-4,
-41,
-127,
-147,
-18,
-8,
-255,
-62,
-175,
-46,
-79,
-138,
-88,
-98,
-26,
-41,
-219,
-39,
-58,
-100,
-157,
-117,
-127,
-124,
-170,
-61,
187,
187,
200,
246,
233,
78,
179,
229,
210,
240,
215,
249,
51,
45,
215,
193,
73,
31,
182,
188,
204,
32,
168,
114,
135,
174,
163,
154,
22,
205,
81,
124,
168,
153,
47,
147,
24,
228,
142,
234,
8,
67,
180,
225,
4,
177,
227,
197,
124,
88,
177,
12,
125,
69,
227,
203,
148,
90,
28,
220,
207,
236,
-146,
-197,
-224,
-13,
-225,
-36,
-128,
-151,
-200,
-69,
-195,
-2,
-232,
-91,
-37,
-71,
-100,
-8,
-75,
-90,
-131,
-93,
-142,
-206,
-197,
-55,
-181,
-220,
-159,
-2,
-15,
-227,
-32,
-252,
-30,
-160,
-112,
-3,
-188,
-65,
-246,
-249,
-227,
-204,
-152,
-42,
-45,
-187,
-72,
-42,
-188,
-27,
-100,
-239,
-243,
-99,
-64,
-35,
-22,
-233,
-160,
-16,
-169,
91,
83,
215,
11,
61,
17,
181,
88,
40,
90,
88,
164,
192,
122,
153,
124,
175,
9,
53,
194,
55,
123,
232,
205,
97,
0,
164,
228,
202,
146,
23,
209,
64,
163,
148,
74,
204,
216,
196,
75,
98,
119,
32,
184,
88,
139,
132,
112,
152,
246,
35,
238,
133,
210,
158,
23,
224,
88,
167,
52,
119,
251,
-107,
-145,
-131,
-48,
-96,
-210,
-216,
-22,
-137,
-54,
-24,
-68,
-114,
-161,
-5,
-214,
-32,
-99,
-180,
-185,
-56,
-216,
-36,
-197,
-57,
-233,
-217,
-22,
-186,
-236,
-28,
-88,
-79,
-190,
-36,
-109,
-109,
-196,
-158,
-184,
-63,
-9,
-256,
-161,
-113,
-74,
-3,
-173,
-141,
-241,
-37,
-124,
-184,
-9,
-69,
-243,
-96,
-236,
-46,
-28,
-68,
-67,
-185,
246,
137,
210,
171,
-1,
236,
248,
154,
3,
51,
85,
163,
219,
164,
222,
48,
156,
210,
164,
237,
238,
144,
198,
153,
242,
199,
39,
179,
58,
220,
198,
32,
106,
230,
184,
142,
127,
176,
93,
139,
147,
190,
156,
166,
56,
242,
32,
173,
142,
136,
94,
91,
227,
199,
32,
89,
56,
180,
154,
190,
171,
120,
-203,
-25,
-226,
-77,
-88,
-208,
-212,
-3,
-54,
-57,
-216,
-123,
-27,
-47,
-45,
-226,
-138,
-64,
-256,
-4,
-223,
-97,
-175,
-123,
-181,
-157,
-7,
-17,
-104,
-215,
-104,
-101,
-108,
-74,
-141,
-91,
-175,
-81,
-65,
-151,
-239,
-251,
-201,
-62,
-26,
-194,
-99,
-30,
-133,
-30,
-5,
-82,
-38,
-67,
-182,
-69,
-119,
-102,
-204,
-44,
-232,
-3,
-241,
174,
23,
84,
56,
131,
68,
178,
183,
69,
39,
191,
166,
191,
8,
29,
34,
243,
20,
26,
75,
204,
67,
10,
105,
42,
108,
254,
43,
4,
147,
247,
206,
181,
98,
210,
84,
145,
209,
109,
47,
157,
240,
230,
31,
58,
166,
238,
62,
20,
175,
25,
229,
198,
44,
220,
227,
140,
98,
74,
226,
180,
205,
-117,
-71,
-98,
-168,
-75,
-245,
-195,
-119,
-136,
-72,
-19,
-130,
-21,
-220,
-26,
-66,
-47,
-61,
-152,
-142,
-3,
-147,
-5,
-256,
-252,
-105,
-96,
-115,
-154,
-61,
-30,
-36,
-34,
-45,
-209,
-88,
-52,
-236,
-61,
-196,
-72,
-24,
-10,
-22,
-179,
-10,
-26,
-185,
-11,
-4,
-45,
-203,
-148,
-54,
-112,
-182,
-112,
-109,
-112,
-92,
-158,
-87,
-15
);

----------------------------------------------------------------------------------
BEGIN
----------------------------------------------------------------------------------

  PROCESS(aclk) BEGIN
    IF rising_edge(aclk) THEN
      IF s_axis_data_tvalid = '1' THEN
        IF NOT (STD_LOGIC_VECTOR(TO_SIGNED(C_FIR_IN(cnt_fir_in),s_axis_data_tdata'LENGTH)) = s_axis_data_tdata) THEN
          REPORT LF & "----------------------------------------------------------------------------------" & LF &
                 "ERROR: Mismatch of input data! Expected data " &
                 INTEGER'image(C_FIR_IN(cnt_fir_in)) &
                 ", actual data " &
                 INTEGER'image(TO_INTEGER(SIGNED(s_axis_data_tdata))) &
                 LF & "----------------------------------------------------------------------------------" & LF
          SEVERITY ERROR;
        END IF;
        cnt_fir_in <= cnt_fir_in + 1;
      END IF;
    END IF;
  END PROCESS;


  --------------------------------------------------------------------------------

  PROCESS(aclk) BEGIN
    IF rising_edge(aclk) THEN
      s_axis_data_tvalid_i  <= s_axis_data_tvalid;
      s_axis_data_tvalid_ii <= s_axis_data_tvalid_i;
      m_axis_data_tvalid    <= s_axis_data_tvalid_ii;

      IF s_axis_data_tvalid_ii = '1' THEN

        IF cnt_fir_out = 999 THEN
          cnt_fir_out <= 0;
        ELSE
          cnt_fir_out <= cnt_fir_out + 1;
        END IF;

        m_axis_data_tdata <= STD_LOGIC_VECTOR(TO_SIGNED(C_FIR_RESPONSE(cnt_fir_out),m_axis_data_tdata'LENGTH));

      END IF;


    END IF;
  END PROCESS;

  s_axis_data_tready <= '1';

----------------------------------------------------------------------------------
END structural;
----------------------------------------------------------------------------------
