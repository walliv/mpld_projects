----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
----------------------------------------------------------------------------------
ENTITY RP_top IS
  PORT(
    BTN             : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
    SW              : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
    LED             : OUT STD_LOGIC_VECTOR (7 DOWNTO 0) := (others => '0')
  );
END RP_top;
----------------------------------------------------------------------------------
ARCHITECTURE Structural OF RP_top IS
----------------------------------------------------------------------------------



----------------------------------------------------------------------------------
BEGIN
----------------------------------------------------------------------------------

    simple_adder_i : entity work.simple_adder
    generic map(
        WIDTH => 4
    )
    port map(
        A => SW,
        B => BTN,
        Y => LED(3 downto 0),
        C => LED(4),
        Z => LED(7)
    );

----------------------------------------------------------------------------------
END Structural;
----------------------------------------------------------------------------------
